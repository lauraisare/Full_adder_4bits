library verilog;
use verilog.vl_types.all;
entity formula_vlg_vec_tst is
end formula_vlg_vec_tst;
